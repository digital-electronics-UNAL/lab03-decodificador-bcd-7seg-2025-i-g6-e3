`include "sum/sum8b.v"

module sumyrest(
    input [7:0] A,
    input [7:0] B,
    input Sel,
    output CO,
    output [7:0] S0
); // parentesis vacio porque no tiene entradas ni salidas


    wire X0, X1, X2, X3, X4, X5, X6, X7;
    wire [7:0] B2;

    xor(X0,Sel,B[0]);
    xor(X1,Sel,B[1]);
    xor(X2,Sel,B[2]);
    xor(X3,Sel,B[3]);
    xor(X4,Sel,B[4]);
    xor(X5,Sel,B[5]);
    xor(X6,Sel,B[6]);
    xor(X7,Sel,B[7]);

    assign B2[0] = X0;
    assign B2[1] = X1;
    assign B2[2] = X2;
    assign B2[3] = X3;
    assign B2[4] = X4;
    assign B2[5] = X5;
    assign B2[6] = X6;
    assign B2[7] = X7;
    
    sum8b S1 ( 
        .A(A),.B(B2),.Ci(Sel),.CO(CO),.S0(S0)
    ); 

endmodule